module cache#(parameter BITS_DATA = 32, BITS_ADDRESS = 32, ASSOCIATIVITY = 2)
(
    
);

endmodule