module mod_unit
(
    input logic in, mod,
    output logic out
);


endmodule